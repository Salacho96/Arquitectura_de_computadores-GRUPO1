library verilog;
use verilog.vl_types.all;
entity FLIP_FLOP_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end FLIP_FLOP_vlg_check_tst;
