library verilog;
use verilog.vl_types.all;
entity FLIP_FLOP_vlg_vec_tst is
end FLIP_FLOP_vlg_vec_tst;
